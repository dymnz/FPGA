module Multiplxer