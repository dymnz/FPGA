module DFF_N module counter #(parameter WIDTH = 8) (D, CLK, RST, Q)


endmodule